library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is

-- CONSTANTES NUMERICAS

constant tamBus:		integer := 3;

end constants;
